LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY BCDDisplay IS
	PORT (
		V : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		HEX01 : OUT STD_LOGIC_VECTOR(0 TO 6);
		HEX00 : OUT STD_LOGIC_VECTOR(0 TO 6)
	);
END ENTITY;

ARCHITECTURE behave OF BCDDisplay IS
	SIGNAL digit1, digit0 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	COMPONENT BCD IS
		PORT (
			c : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			HEXn : OUT STD_LOGIC_VECTOR(0 TO 6)
		);
	END COMPONENT;
BEGIN
	digit1 <= STD_LOGIC_VECTOR(unsigned(V) / 10)(3 DOWNTO 0);
	digit0 <= STD_LOGIC_VECTOR(unsigned(V) MOD 10)(3 DOWNTO 0);
	HEXn1 : BCD PORT MAP(c => digit1, HEXn => HEX01);
	HEXn0 : BCD PORT MAP(c => digit0, HEXn => HEX00);
END ARCHITECTURE;