LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY AddSub IS
    PORT (
        SIGNAL A, B : IN STD_LOGIC_VECTOR(8 DOWNTO 0);
        SIGNAL sel : IN STD_LOGIC;
        SIGNAL C : OUT STD_LOGIC_VECTOR(8 DOWNTO 0)
    );
END AddSub;

ARCHITECTURE arch OF AddSub IS
BEGIN
C <= STD_LOGIC_VECTOR(UNSIGNED(A) + UNSIGNED(B)) WHEN sel = '0' ELSE
        STD_LOGIC_VECTOR(UNSIGNED(A) - UNSIGNED(B));
END ARCHITECTURE;